BZh91AY&SY�L� 
߀Px����߰?���PX�32
P54I�D��� ���  昙2h�`��` ���DD�T2z�
xI��@ &��bdɣ	�bi�L#0	"H0#I���i��@ 6�ҁ@*��$3����hl@�>���ZK�£�.a��F�\�=~$���q�u��&���⤩��F%�vF[h"��)E8 ��u��O�A��7����$���oqE��v7�o��`�F���b�&L�a�Z���L|�c"�y]�1���l��}� ڿ���L�TVk�3�m	(YZd�z�f��[�1jN��*���!�! �ƥ�8�N�	����䟭��P�N5�gu�[��!���a�!�`�P�������@qp�"a��d��2��r��&�L~�����1�h��h},��:�20AH�;�4���=��ғ~Q$���[�琇�yA;�i�(�pL�P�L9#����"8�]��?0@ʺ��T�͜�N|~���QR�e�T0c�5�^�I�Ñ�H:Q�	���I�X���,1���Q<
���bH�Ɲcn���j]	1�+��d�9���AV����-n�"3�,�ٜ� Hi�,0�+d�2���[	��X�o�Ó_-P<�a]�(9�J��m�7n��!��<�P�0��5��i�v[:��r���uc���&L�
BLQID)ש�7�m(͛O�v�W��Q
`�S;B�9-�My��R�/����V�̝@�G-D��e�Ax���&/݊Sb��\0̃`�rԉ��w$S�	�́0